module XOR2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule

module AND2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule

module AO22X1 (IN1,IN2,IN3,IN4,Q);
	input IN1,IN2,IN3,IN4
	output Q
endmodule
